/*
	Marina Ring, mring@hmc.edu, 10/28/24
	Module to test the AES controller module
	
*/

module testbench_aes_controller();
	logic [127:0] key;
	logic clk, load;
	logic sben, sben_expected, sren, sren_expected, mcen, mcen_expected, outen, outen_expected, done, done_expected;
	logic [127:0] roundkey, roundkey_expected;

	logic [31:0] vectornum, errors;
	logic [261:0] testvectors[10000:0];
	
	aes_controller controller(clk, key, sben, sren, mcen, outen, done, roundkey);
	
	always 
		begin
			clk = 1; #5; clk = 0; #5;
		end
	
	initial 
		begin
			$readmemh("aes_controller_tv.txt", testvectors); // readmemh ensures that we can write aes_controller in hexadecimal!!!
			vectornum = 0; errors = 0;
			load = 0; #22; load = 1;
		end
	
	always @(posedge clk)
		begin
			#1; {load, key, sben_expected, sren_expected, mcen_expected, outen_expected, done_expected, roundkey_expected} = testvectors[vectornum];
		end
		
	always @(negedge clk)
		if (load) begin // skip during reset
			if (sben_expected != sben || sren_expected != sren || mcen_expected != mcen || outen_expected != outen || done_expected != done) begin // check result
				$display("Error: input = %b", {load, key});
				$display(" outputs = %b (%b expected)", {sben, sren, mcen, outen, done}, {sben_expected, sren_expected, mcen_expected, outen_expected, done_expected});
				errors = errors + 1;
			end
			if (roundkey_expected != roundkey) begin
				$display("Error: input = %h", {load, key});
				$display(" outputs = %h (%h expected)", {roundkey}, {roundkey_expected});
				errors = errors + 1;
			end
			vectornum = vectornum + 1;
			if (testvectors[vectornum] === 262'hx) begin
				$display("%d tests completed with %d errors", vectornum, errors);
				$stop;
			end
		end
endmodule
