/*
	Marina Ring, mring@g.hmc.edu, 10/27/2024
	Module that will call rotation of bytes within each word
*/

